`timescale 1ns / 1ps

module datapath(

    );
endmodule
